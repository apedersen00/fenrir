package conv_pkg;

    // CONVOLUTION PARAMETERS
    parameter int DEFAULT_KERNEL_SIZE = 3;
    parameter int DEFAULT_IN_CHANNELS = 2;
    parameter int DEFAULT_OUT_CHANNELS = 2;
    parameter int DEFAULT_IMG_HEIGHT = 8;
    parameter int DEFAULT_IMG_WIDTH = 8;

    // MEMORY PARMETERS 
    parameter int DEFAULT_BITS_PER_KERNEL_WEIGHT = 6;
    parameter int DEFAULT_BITS_PER_COORDINATE = 4;
    

endpackage