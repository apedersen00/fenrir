library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.conv_pool_pkg.all;

entity conv_pool is
    generic(
        CHANNELS_IN : integer := 1;
        CHANNELS_OUT : integer := 1;
        BITS_PER_NEURON : integer := 6;
        BITS_PER_WEIGHT : integer := 6;
        IMG_WIDTH : integer := 32;
        IMG_HEIGHT : integer := 32;
        BITS_PER_COORD : integer := 8
    );
    port(
        -- Standard ports needed for digital components
        clk : in std_logic;
        rst_i : in std_logic;
        enable_i : in std_logic;

        -- Control signals
        timestep_i : in std_logic;

        -- Event signals
        event_fifo_empty_i : in std_logic;
        event_fifo_bus_i : in std_logic_vector(2 * BITS_PER_COORD + CHANNELS_IN - 1 downto 0);
        event_fifo_read_o : out std_logic;

        -- pragma translate_off
        debug_main_state : out main_state_et;
        debug_next_state : out main_state_et;
        debug_last_state : out main_state_et;
        
        debug_timestep_pending : out std_logic;
        debug_current_event : out event_tensor_t;
        debug_event_valid : out std_logic;
        debug_read_cycle : out integer; -- NEW: Debug signal to show which cycle we're in
        debug_main_state_vec, debug_next_state_vec, debug_last_state_vec : out std_logic_vector(2 downto 0)
        -- pragma translate_on
    );
end entity conv_pool;

architecture rtl of conv_pool is

    signal main_state, main_next_state, main_last_state : main_state_et := IDLE;
    signal timestep_pending : std_logic := '0';
    
    signal current_event : event_tensor_t := (
        x_coord => 0,
        y_coord => 0,
        channel => 0
    );
    signal event_valid : std_logic := '0';
    
    -- NEW: Counter to track cycles within READ_REQUEST state
    signal read_cycle_counter : integer range 1 to 2 := 1;

begin

    -- UPDATED: Read request logic for 2-cycle protocol
    event_fifo_read_o <= '1' when (main_state = READ_REQUEST and read_cycle_counter = 1) else '0';

    state_register_update : process (clk, rst_i)
    begin
        if rising_edge(clk) then
            if rst_i = '1' then
                main_state <= RESET;
            else
                main_state <= main_next_state;
            end if;
        end if;
    end process state_register_update;

    update_last_state : process (clk, rst_i)
    begin
        if rising_edge(clk) then
            if rst_i = '1' then
                main_last_state <= IDLE;
            elsif main_state /= PAUSE then
                main_last_state <= main_state;
            end if;
        end if;
    end process update_last_state;

    -- UPDATED: State machine with 2-cycle READ_REQUEST handling
    state_machine_control : process (all)
    begin
        main_next_state <= main_state; -- Default: stay in current state

        if enable_i = '0' then
            main_next_state <= PAUSE;
        else
            case main_state is
            when IDLE =>
                -- Priority 1: Check timestep
                if timestep_pending = '1' then
                    main_next_state <= POOL;
                -- Priority 2: Check FIFO 
                elsif event_fifo_empty_i = '0' then
                    main_next_state <= READ_REQUEST;
                end if;
                
            when READ_REQUEST =>
                -- Stay in READ_REQUEST for 2 cycles, then go to EVENT_CONV
                if read_cycle_counter = 2 then
                    main_next_state <= EVENT_CONV;
                end if;
                
            when EVENT_CONV => 
                -- Process event, then back to IDLE
                main_next_state <= IDLE;
                
            when PAUSE => 
                main_next_state <= main_last_state;
                
            when POOL =>
                -- Pool processing, then back to IDLE
                main_next_state <= IDLE;
                
            when CONFIG =>
                main_next_state <= IDLE;
                
            when RESET => 
                main_next_state <= IDLE;
            end case;
        end if;
    end process state_machine_control;

    timestep_buffer : process (clk, rst_i)
    begin
        if rising_edge(clk) then
            if rst_i = '1' then 
                timestep_pending <= '0';
            else
                if timestep_i = '1' then
                    timestep_pending <= '1';
                elsif main_state = POOL then
                    timestep_pending <= '0';
                end if;
            end if;
        end if;
    end process timestep_buffer;

    -- NEW: Read cycle counter management
    read_cycle_management : process (clk, rst_i)
    begin
        if rising_edge(clk) then
            if rst_i = '1' then
                read_cycle_counter <= 1;
            else
                if main_state = READ_REQUEST then
                    if read_cycle_counter < 2 then
                        read_cycle_counter <= read_cycle_counter + 1;
                    end if;
                else
                    read_cycle_counter <= 1; -- Reset counter when leaving READ_REQUEST
                end if;
            end if;
        end if;
    end process read_cycle_management;

    -- UPDATED: Event capture process with proper timing
    event_capture : process (clk, rst_i)
    begin
        if rising_edge(clk) then
            if rst_i = '1' then 
                current_event <= (x_coord => 0, y_coord => 0, channel => 0);
                event_valid <= '0';
            else
                -- Capture event on cycle 2 of READ_REQUEST (when FIFO data is valid)
                if main_state = READ_REQUEST and read_cycle_counter = 2 then
                    current_event <= bus_to_event_tensor(
                        event_fifo_bus_i,
                        BITS_PER_COORD,
                        CHANNELS_IN
                    );
                    event_valid <= '1';
                end if;
                
                -- Clear when returning to IDLE
                if main_state = EVENT_CONV and main_next_state = IDLE then
                    event_valid <= '0';
                end if;
            end if;
        end if;
    end process event_capture;

    -- pragma translate_off
    debug_main_state <= main_state;
    debug_next_state <= main_next_state;
    debug_last_state <= main_last_state;
    debug_timestep_pending <= timestep_pending;
    debug_current_event <= current_event;
    debug_event_valid <= event_valid;
    debug_read_cycle <= read_cycle_counter; -- NEW: Debug the cycle counter
    debug_main_state_vec <= state_to_slv(main_state);
    debug_next_state_vec <= state_to_slv(main_next_state);
    debug_last_state_vec <= state_to_slv(main_last_state);
    -- pragma translate_on

end architecture rtl;