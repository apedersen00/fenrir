import snn_interfaces_pkg::*;

module tb_conv_multichannel;

    localparam int COORD_BITS = 3; // address space 0-7
    localparam int IN_CHANNELS = 2;
    localparam int OUT_CHANNELS = 2;
    localparam int KERNEL_SIZE = 3;
    localparam int IMG_WIDTH = 8;
    localparam int IMG_HEIGHT = 8;

    

endmodule