library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_convolution_layer is
end entity tb_convolution_layer;

