package conv_pkg;

    typedef enum logic{
        MUX_CONVOLUTION,
        MUX_POOLING
    } arbiter_mode_t;

endpackage